`include "params.sv"
`include "mem.sv"
`include "mem_interface.sv"
`include "mem_trans.sv"
`include "mem_monitor.sv" 
`include "mem_scb.sv"
`include "mem_driver.sv" 
`include "driver_v2.sv"
`include "test.sv"
`include "mem_tb_top.sv"